`defeine IDLE 0
`define START 1
`define TX    2
`define RX 	  3
`define STOP  4
`define WAIT  5


module i2c(clk,csn,addr,wrn,d_in,rdn,d_out,sda,scl,i2c_clk,
	pulse_counbt,bit_count,curr_state,next_state);

	
endmodule